module onebitshift_64(in64, out64);
	input [63:0] in64;
	output [63:0] out64;

	assign out64[0] = 1'b0;
	assign out64[1] = in64[0];
	assign out64[2] = in64[1];
	assign out64[3] = in64[2];
	assign out64[4] = in64[3];
	assign out64[5] = in64[4];
	assign out64[6] = in64[5];
	assign out64[7] = in64[6];
	assign out64[8] = in64[7];
	assign out64[9] = in64[8];
	assign out64[10] = in64[9];
	assign out64[11] = in64[10];
	assign out64[12] = in64[11];
	assign out64[13] = in64[12];
	assign out64[14] = in64[13];
	assign out64[15] = in64[14];
	assign out64[16] = in64[15];
	assign out64[17] = in64[16];
	assign out64[18] = in64[17];
	assign out64[19] = in64[18];
	assign out64[20] = in64[19];
	assign out64[21] = in64[20];
	assign out64[22] = in64[21];
	assign out64[23] = in64[22];
	assign out64[24] = in64[23];
	assign out64[25] = in64[24];
	assign out64[26] = in64[25];
	assign out64[27] = in64[26];
	assign out64[28] = in64[27];
	assign out64[29] = in64[28];
	assign out64[30] = in64[29];
	assign out64[31] = in64[30];
	assign out64[32] = in64[31];
	assign out64[33] = in64[32];
	assign out64[34] = in64[33];
	assign out64[35] = in64[34];
	assign out64[36] = in64[35];
	assign out64[37] = in64[36];
	assign out64[38] = in64[37];
	assign out64[39] = in64[38];
	assign out64[40] = in64[39];
	assign out64[41] = in64[40];
	assign out64[42] = in64[41];
	assign out64[43] = in64[42];
	assign out64[44] = in64[43];
	assign out64[45] = in64[44];
	assign out64[46] = in64[45];
	assign out64[47] = in64[46];
	assign out64[48] = in64[47];
	assign out64[49] = in64[48];
	assign out64[50] = in64[49];
	assign out64[51] = in64[50];
	assign out64[52] = in64[51];
	assign out64[53] = in64[52];
	assign out64[54] = in64[53];
	assign out64[55] = in64[54];
	assign out64[56] = in64[55];
	assign out64[57] = in64[56];
	assign out64[58] = in64[57];
	assign out64[59] = in64[58];
	assign out64[60] = in64[59];
	assign out64[61] = in64[60];
	assign out64[62] = in64[61];
	assign out64[63] = in64[62];

endmodule