module twos_complement_flipper32(x, xout);
	input [31:0] x;
	output [31:0] xout;
	not notter0(xout[0], x[0]);
	not notter1(xout[1], x[1]);
	not notter2(xout[2], x[2]);
	not notter3(xout[3], x[3]);
	not notter4(xout[4], x[4]);
	not notter5(xout[5], x[5]);
	not notter6(xout[6], x[6]);
	not notter7(xout[7], x[7]);
	not notter8(xout[8], x[8]);
	not notter9(xout[9], x[9]);
	not notter10(xout[10], x[10]);
	not notter11(xout[11], x[11]);
	not notter12(xout[12], x[12]);
	not notter13(xout[13], x[13]);
	not notter14(xout[14], x[14]);
	not notter15(xout[15], x[15]);
	not notter16(xout[16], x[16]);
	not notter17(xout[17], x[17]);
	not notter18(xout[18], x[18]);
	not notter19(xout[19], x[19]);
	not notter20(xout[20], x[20]);
	not notter21(xout[21], x[21]);
	not notter22(xout[22], x[22]);
	not notter23(xout[23], x[23]);
	not notter24(xout[24], x[24]);
	not notter25(xout[25], x[25]);
	not notter26(xout[26], x[26]);
	not notter27(xout[27], x[27]);
	not notter28(xout[28], x[28]);
	not notter29(xout[29], x[29]);
	not notter30(xout[30], x[30]);
	not notter31(xout[31], x[31]);


endmodule