module onebitshift_32(in32, out32);
	input [31:0] in32;
	output [31:0] out32;
	
	assign out32[0] = 0;
	assign out32[1] = in32[0];
	assign out32[2] = in32[1];
	assign out32[3] = in32[2];
	assign out32[4] = in32[3];
	assign out32[5] = in32[4];
	assign out32[6] = in32[5];
	assign out32[7] = in32[6];
	assign out32[8] = in32[7];
	assign out32[9] = in32[8];
	assign out32[10] = in32[9];
	assign out32[11] = in32[10];
	assign out32[12] = in32[11];
	assign out32[13] = in32[12];
	assign out32[14] = in32[13];
	assign out32[15] = in32[14];
	assign out32[16] = in32[15];
	assign out32[17] = in32[16];
	assign out32[18] = in32[17];
	assign out32[19] = in32[18];
	assign out32[20] = in32[19];
	assign out32[21] = in32[20];
	assign out32[22] = in32[21];
	assign out32[23] = in32[22];
	assign out32[24] = in32[23];
	assign out32[25] = in32[24];
	assign out32[26] = in32[25];
	assign out32[27] = in32[26];
	assign out32[28] = in32[27];
	assign out32[29] = in32[28];
	assign out32[30] = in32[29];
	assign out32[31] = in32[30];
 
endmodule